Half Adder block
*
vdd 8 0 dc 5v
*for voltage 5v
vin 1 0 dc 0 PULSE(0 5 0 0.1NS 0.1NS 50NS 100NS)
*input 1
vina 2 0 dc 0 PULSE(0 5 0 0.1NS 0.1NS 100NS 200NS)
*input 2
.SUBCKT NAND 1 4 2 3
m1 3 1 2 2 p1
m2 3 4 2 2 p1
m3 3 1 5 0 n1
m4 5 4 0 0 n1
.ENDS NAND
*
X1 1 2 8 3 NAND
X2 1 3 8 5 NAND
X3 3 2 8 6 NAND
X4 5 6 8 7 NAND
X5 3 3 8 4 NAND
* Output 1 node is 7
* Output 2 node is 4
.model p1 PMOS W=10u
.model n1 NMOS W=10u
.tran 0.001Ns 400Ns
*voltage simulation
.control
*
set color0 = white
set color1 = black
set color2 = blue
set color3 = red
set color4 = orange
set color5 = teal
set xbrushwidth=3
run
plot 18+v(7) 12+v(4) v(1) 6+v(2) 
.endc
.end
*EE19BTECH11041
