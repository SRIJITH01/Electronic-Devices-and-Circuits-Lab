Not Gate
*
vdd 3 0 dc 5v
vin 1 0 dc 0v
*for voltage 5v
m1 2 1 3 3 p1
m2 2 1 0 0 n1
*
.model p1 PMOS W=1u
.model n1 NMOS W=10u
.dc vin 0 5 0.01
*voltage simulation
.control
*
set color0 = white
set color1 = black
set color2 = blue
set xbrushwidth=2
run
plot v(2) vs v(1)
.endc
.end
*EE19BTECH11041